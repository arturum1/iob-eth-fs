// general_operation: General operation group
// Core Configuration Macros.
`define IOB_COVERAGE_ANALYZE_VERSION 16'h0081
