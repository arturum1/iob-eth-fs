// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_RAM_TDP_HEXFILE "none"
`define IOB_RAM_TDP_ADDR_W 6
`define IOB_RAM_TDP_DATA_W 8
`define IOB_RAM_TDP_MEM_NO_READ_ON_WRITE 1
// Core Configuration Macros.
`define IOB_RAM_TDP_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_RAM_TDP_MEM_INIT_FILE_INT HEXFILE
