// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_CTLS_W 21
`define IOB_CTLS_MODE 0
`define IOB_CTLS_SYMBOL 0
// Core Configuration Macros.
`define IOB_CTLS_VERSION 16'h0081
