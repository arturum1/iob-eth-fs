// general_operation: General operation group
// Core Configuration Macros.
`define IOB_ETH_RX_VERSION 16'h0081
