// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXI_INTERCONNECT_ID_WIDTH 8
`define IOB_AXI_INTERCONNECT_DATA_WIDTH 32
`define IOB_AXI_INTERCONNECT_ADDR_WIDTH 32
`define IOB_AXI_INTERCONNECT_M_ADDR_WIDTH 32
`define IOB_AXI_INTERCONNECT_S_COUNT 4
`define IOB_AXI_INTERCONNECT_M_COUNT 4
// Core Configuration Macros.
`define IOB_AXI_INTERCONNECT_VERSION 16'h0081
