// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_GRAY_COUNTER_W 1
// Core Configuration Macros.
`define IOB_GRAY_COUNTER_VERSION 16'h0081
