// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXISTREAM_IN_DATA_W 32
`define IOB_AXISTREAM_IN_ADDR_W 5
`define IOB_AXISTREAM_IN_TDATA_W 8
`define IOB_AXISTREAM_IN_FIFO_ADDR_W 4
// Core Configuration Macros.
`define IOB_AXISTREAM_IN_VERSION 16'h0081
