// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_SYNC_REG_A_DATA_W 1
`define IOB_SYNC_REG_A_RST_VAL {DATA_W{1'b0}}
// Core Configuration Macros.
`define IOB_SYNC_REG_A_VERSION 16'h0001
