// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_AXIS_S_AXI_M_AXI_ADDR_W 1
`define IOB_AXIS_S_AXI_M_AXI_LEN_W 8
`define IOB_AXIS_S_AXI_M_AXI_DATA_W 32
`define IOB_AXIS_S_AXI_M_AXI_ID_W 1
`define IOB_AXIS_S_AXI_M_WLEN_W 1
`define IOB_AXIS_S_AXI_M_RLEN_W 1
// Core Configuration Macros.
`define IOB_AXIS_S_AXI_M_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_AXIS_S_AXI_M_WRITE_HEXFILE "none"
`define IOB_AXIS_S_AXI_M_READ_HEXFILE "none"
