// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_FIFO2AXIS_DATA_W 1
`define IOB_FIFO2AXIS_AXIS_LEN_W 1
// Core Configuration Macros.
`define IOB_FIFO2AXIS_VERSION 16'h0081
