// general_operation: General operation group
// Core Configuration Macros.
`define TB_PBUS_SPLIT_VERSION 16'h0081
