// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_ETH_CSRS_DATA_W 32
`define IOB_ETH_CSRS_AXI_ID_W 1
`define IOB_ETH_CSRS_AXI_ADDR_W 24
`define IOB_ETH_CSRS_AXI_DATA_W 32
`define IOB_ETH_CSRS_AXI_LEN_W 4
`define IOB_ETH_CSRS_PHY_RST_CNT 20'hFFFFF
`define IOB_ETH_CSRS_BD_NUM_LOG2 7
`define IOB_ETH_CSRS_BUFFER_W 11
// Core Configuration Macros.
`define IOB_ETH_CSRS_PREAMBLE 8'h55
`define IOB_ETH_CSRS_PREAMBLE_LEN 7
`define IOB_ETH_CSRS_SFD 8'hD5
`define IOB_ETH_CSRS_MAC_ADDR_LEN 6
`define IOB_ETH_CSRS_MODER_ADDR 0
`define IOB_ETH_CSRS_MODER_W 32
`define IOB_ETH_CSRS_INT_SOURCE_ADDR 4
`define IOB_ETH_CSRS_INT_SOURCE_W 32
`define IOB_ETH_CSRS_INT_MASK_ADDR 8
`define IOB_ETH_CSRS_INT_MASK_W 32
`define IOB_ETH_CSRS_IPGT_ADDR 12
`define IOB_ETH_CSRS_IPGT_W 32
`define IOB_ETH_CSRS_IPGR1_ADDR 16
`define IOB_ETH_CSRS_IPGR1_W 32
`define IOB_ETH_CSRS_IPGR2_ADDR 20
`define IOB_ETH_CSRS_IPGR2_W 32
`define IOB_ETH_CSRS_PACKETLEN_ADDR 24
`define IOB_ETH_CSRS_PACKETLEN_W 32
`define IOB_ETH_CSRS_COLLCONF_ADDR 28
`define IOB_ETH_CSRS_COLLCONF_W 32
`define IOB_ETH_CSRS_TX_BD_NUM_ADDR 32
`define IOB_ETH_CSRS_TX_BD_NUM_W 32
`define IOB_ETH_CSRS_CTRLMODER_ADDR 36
`define IOB_ETH_CSRS_CTRLMODER_W 32
`define IOB_ETH_CSRS_MIIMODER_ADDR 40
`define IOB_ETH_CSRS_MIIMODER_W 32
`define IOB_ETH_CSRS_MIICOMMAND_ADDR 44
`define IOB_ETH_CSRS_MIICOMMAND_W 32
`define IOB_ETH_CSRS_MIIADDRESS_ADDR 48
`define IOB_ETH_CSRS_MIIADDRESS_W 32
`define IOB_ETH_CSRS_MIITX_DATA_ADDR 52
`define IOB_ETH_CSRS_MIITX_DATA_W 32
`define IOB_ETH_CSRS_MIIRX_DATA_ADDR 56
`define IOB_ETH_CSRS_MIIRX_DATA_W 32
`define IOB_ETH_CSRS_MIISTATUS_ADDR 60
`define IOB_ETH_CSRS_MIISTATUS_W 32
`define IOB_ETH_CSRS_MAC_ADDR0_ADDR 64
`define IOB_ETH_CSRS_MAC_ADDR0_W 32
`define IOB_ETH_CSRS_MAC_ADDR1_ADDR 68
`define IOB_ETH_CSRS_MAC_ADDR1_W 32
`define IOB_ETH_CSRS_ETH_HASH0_ADR_ADDR 72
`define IOB_ETH_CSRS_ETH_HASH0_ADR_W 32
`define IOB_ETH_CSRS_ETH_HASH1_ADR_ADDR 76
`define IOB_ETH_CSRS_ETH_HASH1_ADR_W 32
`define IOB_ETH_CSRS_ETH_TXCTRL_ADDR 80
`define IOB_ETH_CSRS_ETH_TXCTRL_W 32
`define IOB_ETH_CSRS_TX_BD_CNT_ADDR 84
`define IOB_ETH_CSRS_TX_BD_CNT_W 8
`define IOB_ETH_CSRS_RX_BD_CNT_ADDR 88
`define IOB_ETH_CSRS_RX_BD_CNT_W 8
`define IOB_ETH_CSRS_TX_WORD_CNT_ADDR 92
`define IOB_ETH_CSRS_TX_WORD_CNT_W 32
`define IOB_ETH_CSRS_RX_WORD_CNT_ADDR 96
`define IOB_ETH_CSRS_RX_WORD_CNT_W 32
`define IOB_ETH_CSRS_RX_NBYTES_ADDR 100
`define IOB_ETH_CSRS_RX_NBYTES_W 32
`define IOB_ETH_CSRS_FRAME_WORD_ADDR 104
`define IOB_ETH_CSRS_FRAME_WORD_W 8
`define IOB_ETH_CSRS_PHY_RST_VAL_ADDR 108
`define IOB_ETH_CSRS_PHY_RST_VAL_W 8
`define IOB_ETH_CSRS_BD_ADDR 1024
`define IOB_ETH_CSRS_BD_W 32
`define IOB_ETH_CSRS_VERSION_ADDR 2048
`define IOB_ETH_CSRS_VERSION_W 16
`define IOB_ETH_CSRS_VERSION 16'h0001
// Core Derived Parameters. DO NOT CHANGE
`define IOB_ETH_CSRS_ADDR_W 12
