// SPDX-FileCopyrightText: 2026 IObundle, Lda
//
// SPDX-License-Identifier: MIT
//
// Py2HWSW Version 0.81 has generated this code (https://github.com/IObundle/py2hwsw).

`timescale 1ns / 1ps
`include "iob_sync_reg_a_conf.vh"

module iob_sync_reg_a #(
   parameter DATA_W  = `IOB_SYNC_REG_A_DATA_W,
   parameter RST_VAL = `IOB_SYNC_REG_A_RST_VAL
) (
   // clk_en_rst_s: Clock, clock enable and reset
   input                   clk_i,
   input                   arst_i,
   // data_i: Data input
   input      [DATA_W-1:0] iob_sync_reg_data_i,
   // data_o: Data output
   output reg [DATA_W-1:0] iob_sync_reg_data_o
);


   always @(posedge clk_i, posedge arst_i) begin
      if (arst_i) begin
         iob_sync_reg_data_o <= RST_VAL;
      end else begin
         iob_sync_reg_data_o <= iob_sync_reg_data_i;
      end
   end



endmodule
