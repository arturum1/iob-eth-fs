// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_DMA_CSRS_DATA_W 32
`define IOB_DMA_CSRS_AXI_ADDR_W 1
`define IOB_DMA_CSRS_AXI_LEN_W 8
`define IOB_DMA_CSRS_AXI_DATA_W 32
`define IOB_DMA_CSRS_AXI_ID_W 1
`define IOB_DMA_CSRS_WLEN_W 12
`define IOB_DMA_CSRS_RLEN_W 12
// Core Configuration Macros.
`define IOB_DMA_CSRS_W_ADDR_ADDR 0
`define IOB_DMA_CSRS_W_ADDR_W 32
`define IOB_DMA_CSRS_W_LENGTH_ADDR 4
`define IOB_DMA_CSRS_W_LENGTH_W 32
`define IOB_DMA_CSRS_W_BUSY_ADDR 0
`define IOB_DMA_CSRS_W_BUSY_W 8
`define IOB_DMA_CSRS_W_START_ADDR 8
`define IOB_DMA_CSRS_W_START_W 8
`define IOB_DMA_CSRS_W_BURSTLEN_ADDR 10
`define IOB_DMA_CSRS_W_BURSTLEN_W 16
`define IOB_DMA_CSRS_W_BUF_LEVEL_ADDR 4
`define IOB_DMA_CSRS_W_BUF_LEVEL_W 32
`define IOB_DMA_CSRS_R_ADDR_ADDR 12
`define IOB_DMA_CSRS_R_ADDR_W 32
`define IOB_DMA_CSRS_R_LENGTH_ADDR 16
`define IOB_DMA_CSRS_R_LENGTH_W 32
`define IOB_DMA_CSRS_R_START_ADDR 20
`define IOB_DMA_CSRS_R_START_W 8
`define IOB_DMA_CSRS_R_BUSY_ADDR 8
`define IOB_DMA_CSRS_R_BUSY_W 8
`define IOB_DMA_CSRS_R_BURSTLEN_ADDR 22
`define IOB_DMA_CSRS_R_BURSTLEN_W 16
`define IOB_DMA_CSRS_R_BUF_LEVEL_ADDR 12
`define IOB_DMA_CSRS_R_BUF_LEVEL_W 32
`define IOB_DMA_CSRS_VERSION_ADDR 16
`define IOB_DMA_CSRS_VERSION_W 16
`define IOB_DMA_CSRS_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_DMA_CSRS_ADDR_W 5
