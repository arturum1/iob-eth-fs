// general_operation: General operation group
// Core Configuration Macros.
`define IOB_LINUX_DEVICE_DRIVERS_VERSION 16'h0081
