// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_MODCNT_DATA_W 21
`define IOB_MODCNT_RST_VAL {DATA_W{1'b0}}
// Core Configuration Macros.
`define IOB_MODCNT_VERSION 16'h0081
