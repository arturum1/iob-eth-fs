// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_ETH_DT_BUFFER_W 11
`define IOB_ETH_DT_BD_ADDR_W 8
// Core Configuration Macros.
`define IOB_ETH_DT_VERSION 16'h0081
// Core Derived Parameters. DO NOT CHANGE
`define IOB_ETH_DT_AXI_ID_W 1
`define IOB_ETH_DT_AXI_LEN_W 8
`define IOB_ETH_DT_AXI_ADDR_W 0
`define IOB_ETH_DT_AXI_DATA_W 32
