// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_GRAY2BIN_DATA_W 4
// Core Configuration Macros.
`define IOB_GRAY2BIN_VERSION 16'h0081
