// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_CLOCK_CLK_PERIOD 10
// Core Configuration Macros.
`define IOB_CLOCK_VERSION 16'h0081
