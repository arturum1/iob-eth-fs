// general_operation: General operation group
// Core Configuration Macros.
`define IOB_ARBITER_VERSION 16'h0081
