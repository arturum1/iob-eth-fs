// general_operation: General operation group
// Core Configuration Macros.
`define IOB_ETH_MII_MANAGEMENT_VERSION 16'h0081
