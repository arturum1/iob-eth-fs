// general_operation: General operation group
// Core Configuration Macros.
`define IOB_RESET_SYNC_VERSION 16'h0081
