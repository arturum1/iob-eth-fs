// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_EDGE_DETECT_EDGE_TYPE "rising"
`define IOB_EDGE_DETECT_OUT_TYPE "step"
// Core Configuration Macros.
`define IOB_EDGE_DETECT_VERSION 16'h0081
